../tme4/adder32b.vhdl