../tme4/alu.vhdl