../tme4/shifter.vhdl